-- 
-- VHDL Architecture proj_master_2025_lib.{$ENTITY_NAME}.struct
--
-- Created at: {$DATE_TIME}
--
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;
{$LIBRARY}


architecture struct of {$ENTITY_NAME} is

   -- Architecture declarations

{$ARCH_DECLARATIONS}

begin
   -- Architecture concurrent statements

{$ARCH_STATEMENTS}

end struct ;