-- VHDL Entity proj_master_2025_lib.{$ENTITY_NAME}.symbol
--
-- Created at: {$DATE_TIME}
--
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

entity {$ENTITY_NAME} is
-- Declarations

end {$ENTITY_NAME} ;