LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;
